  end
  assign rd = ROM[a[31:1]];
endmodule